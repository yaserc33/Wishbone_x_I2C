package i2c_module_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "wb_x_i2c_ref_model.sv"
	`include "i2c_scoreboard.sv"
	`include "i2c_module.sv"
endpackage
